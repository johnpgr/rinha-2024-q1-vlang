module main

@[if debug]
pub fn debug[T](s T) {
	println(s)
}
