module main

fn main() {
	println('Hello World!')
	// init_tables()
	// insert_test_clientes()
}
