module main

@[if debug]
pub fn debug(s string) {
	println(s)
}
